module system

pub const (
	action_farm_define     = 'farmerbot.farmmanager.define'
	action_node_define     = 'farmerbot.nodemanager.define'
	action_power_configure = 'farmerbot.powermanager.configure'
)
