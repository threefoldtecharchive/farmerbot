module system

pub const(
	job_node_find = "farmerbot.nodemanager.find"
)

