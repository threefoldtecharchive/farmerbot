module system

pub const(
	action_node_definition = "farmerbot.node.define"
	action_find_node = "farmerbot.resourcemanager.findnode"
)