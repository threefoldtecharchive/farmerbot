module manager

import freeflowuniverse.baobab.actions
import threefoldtech.farmerbot.system


pub fn data_set(mut db &system.DB, mut action &actions.Action) !{

	// mut node := system.Node{}
	// node.id = action.params.get_u32("id")!
	// node.description = action.params.get_default("description","")!
	// node.farmid = action.params.get_u32("farmid")!
	// node.powermanager = action.params.get("powermanager")!
	// node.powermanager_port = action.params.get_u8("powermanager_port")!
	// db.nodes[node.id]=&node
}