module tasklets



import domain_farmer.actor_capacityplanner
import domain_farmer.actor_powermanager

import domain_tfgrid.actor_notary



// fn (mut tm TaskletManager) action_reboot(mut job &actionrunner.ActionJob)!bool{
