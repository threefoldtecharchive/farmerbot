module system

pub const(
	action_node_define = "farmerbot.nodemanager.define"
)