module actor_notary

const domain="tfgrid"