module system

pub const(
	job_node_find = "farmerbot.nodemanager.find"
	job_power_on = "farmerbot.powermanager.poweron"
)

