module system

pub const(
	job_node_find = "farmerbot.nodemanager.findnode"

	job_power_off = "farmerbot.powermanager.poweroff"
	job_power_on = "farmerbot.powermanager.poweron"
	job_power_periodicwakeup = "farmerbot.powermanager.periodic_wakeup"
	job_power_powermanagement = "farmerbot.powermanager.powermanagement"


)

